LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;
ENTITY ____ IS
	PORT
	( -- put your inputs and outputs here
	   : IN STD_LOGIC;
	   : OUT STD_LOGIC
   )
END ENTITY _________________;

ARCHITECTURE _____ OF  _____  IS

BEGIN

	 ---- enter stuff here
END ARCHITECTURE _____;
